/**
 * Computes the sum of two bits.
 */
CHIP HalfAdder {
    IN a, b;    /* 1-bit inputs */
    OUT sum,    /* Right bit of a + b */
        carry;  /* Left bit of a + b */

    PARTS:
	Xor(a=a, b=b, out=sum);
	And(a=a, b=b, out=carry);
}

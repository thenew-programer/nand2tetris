/**
 * 4-way 16-bit multiplexor:
 * out = a if sel = 00
 *       b if sel = 01
 *       c if sel = 10
 *       d if sel = 11
 */
CHIP Mux4Way16 {
    IN a[16], b[16], c[16], d[16], sel[2];
    OUT out[16];
    
    PARTS:
	Mux16(a=a, b=b, sel=sel[0], out=e);
	Mux16(a=c, b=d, sel=sel[0], out=f);
	Mux16(a=e, b=f, sel=sel[1], out=out);
}

// This file is part of www.nand2tetris.org
// and the book "The Elements of Computing Systems"
// by Nisan and Schocken, MIT Press.
// File name: projects/1/Or.hdl
/**
 * Or gate:
 * if (a or b) out = 1, else out = 0 
 */
CHIP Or {
    IN a, b;
    OUT out;

    PARTS:
	Not(in=a, out=nota);
	Not(in=b, out=notb);
	And(a=nota, b=notb, out=notaAndnotb);
	Not(in=notaAndnotb, out=out);
}
